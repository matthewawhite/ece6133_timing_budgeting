##
## LEF for PtnCells ;
## created by Innovus v17.12-s095_1 on Thu Apr 23 01:11:55 2020
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO Reg_width80
  CLASS BLOCK ;
  FOREIGN Reg_width80 0 0 ;
  ORIGIN 0.0000 0.0000 ;
  SIZE 75.2400 BY 74.1000 ;
  SYMMETRY X Y R90 ;
  PIN input[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 57.4400 0.0700 57.5100 ;
    END
  END input[79]
  PIN input[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 45.0900 0.0700 45.1600 ;
    END
  END input[78]
  PIN input[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 23.4300 74.0300 23.5000 74.1000 ;
    END
  END input[77]
  PIN input[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 50.0300 0.0700 50.1000 ;
    END
  END input[76]
  PIN input[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 18.1100 75.2400 18.1800 ;
    END
  END input[75]
  PIN input[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 70.5500 0.0000 70.6200 0.0700 ;
    END
  END input[74]
  PIN input[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 8.0400 75.2400 8.1100 ;
    END
  END input[73]
  PIN input[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 10.7000 75.2400 10.7700 ;
    END
  END input[72]
  PIN input[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 27.8000 75.2400 27.8700 ;
    END
  END input[71]
  PIN input[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 40.1500 75.2400 40.2200 ;
    END
  END input[70]
  PIN input[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 42.6200 75.2400 42.6900 ;
    END
  END input[69]
  PIN input[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 25.5200 75.2400 25.5900 ;
    END
  END input[68]
  PIN input[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 47.7500 75.2400 47.8200 ;
    END
  END input[67]
  PIN input[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 70.5500 74.0300 70.6200 74.1000 ;
    END
  END input[66]
  PIN input[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 63.3300 74.0300 63.4000 74.1000 ;
    END
  END input[65]
  PIN input[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 51.1700 74.0300 51.2400 74.1000 ;
    END
  END input[64]
  PIN input[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 47.7500 74.0300 47.8200 74.1000 ;
    END
  END input[63]
  PIN input[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.3100 74.0300 52.3800 74.1000 ;
    END
  END input[62]
  PIN input[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.6900 74.0300 33.7600 74.1000 ;
    END
  END input[61]
  PIN input[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 25.3300 74.0300 25.4000 74.1000 ;
    END
  END input[60]
  PIN input[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 40.3400 0.0700 40.4100 ;
    END
  END input[59]
  PIN input[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 37.6800 0.0700 37.7500 ;
    END
  END input[58]
  PIN input[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 30.2700 0.0700 30.3400 ;
    END
  END input[57]
  PIN input[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 53.8300 0.0000 53.9000 0.0700 ;
    END
  END input[56]
  PIN input[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 61.0500 0.0000 61.1200 0.0700 ;
    END
  END input[55]
  PIN input[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 70.5850 0.0000 70.7250 0.1400 ;
    END
  END input[54]
  PIN input[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.4100 0.0000 50.4800 0.0700 ;
    END
  END input[53]
  PIN input[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 12.9800 75.2400 13.0500 ;
    END
  END input[52]
  PIN input[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 37.8700 0.0000 37.9400 0.0700 ;
    END
  END input[51]
  PIN input[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.7900 0.0000 50.8600 0.0700 ;
    END
  END input[50]
  PIN input[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 43.1900 0.0000 43.2600 0.0700 ;
    END
  END input[49]
  PIN input[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 37.6800 75.2400 37.7500 ;
    END
  END input[48]
  PIN input[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 45.4700 74.0300 45.5400 74.1000 ;
    END
  END input[47]
  PIN input[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 62.5700 74.0300 62.6400 74.1000 ;
    END
  END input[46]
  PIN input[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 54.2100 74.0300 54.2800 74.1000 ;
    END
  END input[45]
  PIN input[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 56.8700 74.0300 56.9400 74.1000 ;
    END
  END input[44]
  PIN input[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 43.5700 74.0300 43.6400 74.1000 ;
    END
  END input[43]
  PIN input[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 28.7500 74.0300 28.8200 74.1000 ;
    END
  END input[42]
  PIN input[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 32.1700 74.0300 32.2400 74.1000 ;
    END
  END input[41]
  PIN input[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 42.6200 0.0700 42.6900 ;
    END
  END input[40]
  PIN input[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 34.0700 0.0000 34.1400 0.0700 ;
    END
  END input[39]
  PIN input[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 30.2700 0.0000 30.3400 0.0700 ;
    END
  END input[38]
  PIN input[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.9900 0.0000 28.0600 0.0700 ;
    END
  END input[37]
  PIN input[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 42.4300 0.0000 42.5000 0.0700 ;
    END
  END input[36]
  PIN input[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 45.0900 0.0000 45.1600 0.0700 ;
    END
  END input[35]
  PIN input[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.7700 0.0000 58.8400 0.0700 ;
    END
  END input[34]
  PIN input[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 53.4500 0.0000 53.5200 0.0700 ;
    END
  END input[33]
  PIN input[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 41.6700 0.0000 41.7400 0.0700 ;
    END
  END input[32]
  PIN input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 32.9300 75.2400 33.0000 ;
    END
  END input[31]
  PIN input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 22.8600 75.2400 22.9300 ;
    END
  END input[30]
  PIN input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 35.2100 75.2400 35.2800 ;
    END
  END input[29]
  PIN input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 59.9100 75.2400 59.9800 ;
    END
  END input[28]
  PIN input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 59.8750 75.2400 60.0150 ;
    END
  END input[27]
  PIN input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 47.6200 75.2400 47.7600 ;
    END
  END input[26]
  PIN input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 57.4400 75.2400 57.5100 ;
    END
  END input[25]
  PIN input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 54.0650 73.9600 54.2050 74.1000 ;
    END
  END input[24]
  PIN input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.6900 74.0300 52.7600 74.1000 ;
    END
  END input[23]
  PIN input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 45.3850 73.9600 45.5250 74.1000 ;
    END
  END input[22]
  PIN input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 42.7750 0.1400 42.9150 ;
    END
  END input[21]
  PIN input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.9700 74.0300 36.0400 74.1000 ;
    END
  END input[20]
  PIN input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 32.1700 0.0000 32.2400 0.0700 ;
    END
  END input[19]
  PIN input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 30.2350 0.1400 30.3750 ;
    END
  END input[18]
  PIN input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 22.8600 0.0700 22.9300 ;
    END
  END input[17]
  PIN input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 28.0250 0.0000 28.1650 0.1400 ;
    END
  END input[16]
  PIN input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 18.1100 0.0700 18.1800 ;
    END
  END input[15]
  PIN input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 63.7100 0.0000 63.7800 0.0700 ;
    END
  END input[14]
  PIN input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 49.2700 0.0000 49.3400 0.0700 ;
    END
  END input[13]
  PIN input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 17.9800 75.2400 18.1200 ;
    END
  END input[12]
  PIN input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 15.4500 75.2400 15.5200 ;
    END
  END input[11]
  PIN input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 27.9550 75.2400 28.0950 ;
    END
  END input[10]
  PIN input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 42.7750 75.2400 42.9150 ;
    END
  END input[9]
  PIN input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 47.3950 75.2400 47.7950 ;
    END
  END input[8]
  PIN input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 40.2100 75.2400 40.3500 ;
    END
  END input[7]
  PIN input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 59.1500 74.0300 59.2200 74.1000 ;
    END
  END input[6]
  PIN input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 62.3800 75.2400 62.4500 ;
    END
  END input[5]
  PIN input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.8500 74.0300 64.9200 74.1000 ;
    END
  END input[4]
  PIN input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 40.1500 74.0300 40.2200 74.1000 ;
    END
  END input[3]
  PIN input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 45.8500 74.0300 45.9200 74.1000 ;
    END
  END input[2]
  PIN input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 39.7950 75.2400 40.1950 ;
    END
  END input[1]
  PIN input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.9700 0.0000 36.0400 0.0700 ;
    END
  END input[0]
  PIN output[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 58.9600 0.0700 59.0300 ;
    END
  END output[79]
  PIN output[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 47.7500 0.0700 47.8200 ;
    END
  END output[78]
  PIN output[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 17.5400 74.0300 17.6100 74.1000 ;
    END
  END output[77]
  PIN output[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 57.5950 0.1400 57.7350 ;
    END
  END output[76]
  PIN output[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 24.3800 75.2400 24.4500 ;
    END
  END output[75]
  PIN output[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 60.7850 0.0000 60.9250 0.1400 ;
    END
  END output[74]
  PIN output[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 12.0300 75.2400 12.1000 ;
    END
  END output[73]
  PIN output[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 9.5600 75.2400 9.6300 ;
    END
  END output[72]
  PIN output[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 37.9300 75.2400 38.0700 ;
    END
  END output[71]
  PIN output[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 37.8950 75.2400 38.2950 ;
    END
  END output[70]
  PIN output[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 34.2600 0.0700 34.3300 ;
    END
  END output[69]
  PIN output[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 29.3200 75.2400 29.3900 ;
    END
  END output[68]
  PIN output[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 45.2800 75.2400 45.3500 ;
    END
  END output[67]
  PIN output[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.0100 74.0300 58.0800 74.1000 ;
    END
  END output[66]
  PIN output[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal8 ;
        RECT 53.6550 73.7000 54.0550 74.1000 ;
    END
  END output[65]
  PIN output[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 37.8700 74.0300 37.9400 74.1000 ;
    END
  END output[64]
  PIN output[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 26.4700 74.0300 26.5400 74.1000 ;
    END
  END output[63]
  PIN output[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 47.9050 73.9600 48.0450 74.1000 ;
    END
  END output[62]
  PIN output[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 29.7000 74.0300 29.7700 74.1000 ;
    END
  END output[61]
  PIN output[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 29.4250 73.9600 29.5650 74.1000 ;
    END
  END output[60]
  PIN output[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 40.2100 0.1400 40.3500 ;
    END
  END output[59]
  PIN output[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 35.4000 0.0700 35.4700 ;
    END
  END output[58]
  PIN output[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.2300 0.0000 27.3000 0.0700 ;
    END
  END output[57]
  PIN output[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.3100 0.0000 33.3800 0.0700 ;
    END
  END output[56]
  PIN output[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.4700 0.0000 64.5400 0.0700 ;
    END
  END output[55]
  PIN output[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 55.7300 0.0000 55.8000 0.0700 ;
    END
  END output[54]
  PIN output[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 51.7400 0.0000 51.8100 0.0700 ;
    END
  END output[53]
  PIN output[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 14.5000 75.2400 14.5700 ;
    END
  END output[52]
  PIN output[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.3200 0.0000 48.3900 0.0700 ;
    END
  END output[51]
  PIN output[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 26.8500 75.2400 26.9200 ;
    END
  END output[50]
  PIN output[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal9 ;
        RECT 74.4400 27.0550 75.2400 27.8550 ;
    END
  END output[49]
  PIN output[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT 38.3850 0.0000 38.5250 0.1400 ;
    END
  END output[48]
  PIN output[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.3900 74.0300 58.4600 74.1000 ;
    END
  END output[47]
  PIN output[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 66.5600 74.0300 66.6300 74.1000 ;
    END
  END output[46]
  PIN output[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 54.0200 75.2400 54.0900 ;
    END
  END output[45]
  PIN output[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 56.4900 75.2400 56.5600 ;
    END
  END output[44]
  PIN output[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 45.3400 0.1400 45.4800 ;
    END
  END output[43]
  PIN output[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.0400 74.0300 27.1100 74.1000 ;
    END
  END output[42]
  PIN output[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 42.2400 74.0300 42.3100 74.1000 ;
    END
  END output[41]
  PIN output[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.9900 74.0300 28.0600 74.1000 ;
    END
  END output[40]
  PIN output[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 37.1100 0.0000 37.1800 0.0700 ;
    END
  END output[39]
  PIN output[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 18.6800 0.0000 18.7500 0.0700 ;
    END
  END output[38]
  PIN output[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 16.5900 0.0000 16.6600 0.0700 ;
    END
  END output[37]
  PIN output[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 20.7700 0.0000 20.8400 0.0700 ;
    END
  END output[36]
  PIN output[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT 36.9850 0.0000 37.1250 0.1400 ;
    END
  END output[35]
  PIN output[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 30.6500 0.0000 30.7200 0.0700 ;
    END
  END output[34]
  PIN output[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 51.3600 0.0000 51.4300 0.0700 ;
    END
  END output[33]
  PIN output[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 37.5450 0.0000 37.6850 0.1400 ;
    END
  END output[32]
  PIN output[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 29.0950 75.2400 29.2350 ;
    END
  END output[31]
  PIN output[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 24.5950 75.2400 24.9950 ;
    END
  END output[30]
  PIN output[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 36.7300 75.2400 36.8000 ;
    END
  END output[29]
  PIN output[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 41.6700 75.2400 41.7400 ;
    END
  END output[28]
  PIN output[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 50.2200 75.2400 50.2900 ;
    END
  END output[27]
  PIN output[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 44.1400 75.2400 44.2100 ;
    END
  END output[26]
  PIN output[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 57.5950 75.2400 57.7350 ;
    END
  END output[25]
  PIN output[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 54.0450 75.2400 54.4450 ;
    END
  END output[24]
  PIN output[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 57.4400 74.0300 57.5100 74.1000 ;
    END
  END output[23]
  PIN output[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 41.2900 74.0300 41.3600 74.1000 ;
    END
  END output[22]
  PIN output[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 44.7100 74.0300 44.7800 74.1000 ;
    END
  END output[21]
  PIN output[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 46.6100 75.2400 46.6800 ;
    END
  END output[20]
  PIN output[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 34.1850 0.0000 34.3250 0.1400 ;
    END
  END output[19]
  PIN output[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 39.3900 0.0700 39.4600 ;
    END
  END output[18]
  PIN output[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 37.3600 0.1400 37.5000 ;
    END
  END output[17]
  PIN output[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 0.0000 29.3450 0.4000 29.7450 ;
    END
  END output[16]
  PIN output[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 39.0100 0.0700 39.0800 ;
    END
  END output[15]
  PIN output[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.0900 0.0000 64.1600 0.0700 ;
    END
  END output[14]
  PIN output[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.7000 0.0000 48.7700 0.0700 ;
    END
  END output[13]
  PIN output[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 14.1200 75.2400 14.1900 ;
    END
  END output[12]
  PIN output[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 15.7000 75.2400 15.8400 ;
    END
  END output[11]
  PIN output[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 29.3450 75.2400 29.7450 ;
    END
  END output[10]
  PIN output[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 42.6450 75.2400 43.0450 ;
    END
  END output[9]
  PIN output[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal9 ;
        RECT 74.4400 45.8650 75.2400 46.6650 ;
    END
  END output[8]
  PIN output[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 38.7850 75.2400 38.9250 ;
    END
  END output[7]
  PIN output[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 65.6100 74.0300 65.6800 74.1000 ;
    END
  END output[6]
  PIN output[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 63.9000 75.2400 63.9700 ;
    END
  END output[5]
  PIN output[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 67.5100 74.0300 67.5800 74.1000 ;
    END
  END output[4]
  PIN output[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 37.2650 73.9600 37.4050 74.1000 ;
    END
  END output[3]
  PIN output[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal8 ;
        RECT 47.7750 73.7000 48.1750 74.1000 ;
    END
  END output[2]
  PIN output[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal9 ;
        RECT 74.4400 42.4450 75.2400 43.2450 ;
    END
  END output[1]
  PIN output[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 36.3500 0.0700 36.4200 ;
    END
  END output[0]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 24.9500 0.0700 25.0200 ;
    END
  END enable
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 38.8200 75.2400 38.8900 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 18.8700 0.0700 18.9400 ;
    END
  END reset
  OBS
    LAYER metal10 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal9 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal8 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal7 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal6 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal5 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal4 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal3 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal2 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal1 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
  END
END Reg_width80

END LIBRARY
