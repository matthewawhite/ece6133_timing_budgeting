##
## LEF for PtnCells ;
## created by Innovus v17.12-s095_1 on Wed Apr 22 22:04:46 2020
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AsyncMux_width80
  CLASS BLOCK ;
  FOREIGN AsyncMux_width80 0 0 ;
  ORIGIN 0.0000 0.0000 ;
  SIZE 75.2400 BY 74.1000 ;
  SYMMETRY X Y R90 ;
  PIN input0[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 46.0400 0.0700 46.1100 ;
    END
  END input0[79]
  PIN input0[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 41.1000 0.0700 41.1700 ;
    END
  END input0[78]
  PIN input0[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 43.5700 0.0700 43.6400 ;
    END
  END input0[77]
  PIN input0[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 43.6300 0.1400 43.7700 ;
    END
  END input0[76]
  PIN input0[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 26.2800 75.2400 26.3500 ;
    END
  END input0[75]
  PIN input0[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 50.4250 0.0000 50.5650 0.1400 ;
    END
  END input0[74]
  PIN input0[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 27.4450 75.2400 27.8450 ;
    END
  END input0[73]
  PIN input0[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 28.7500 75.2400 28.8200 ;
    END
  END input0[72]
  PIN input0[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 33.6900 75.2400 33.7600 ;
    END
  END input0[71]
  PIN input0[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 39.7700 75.2400 39.8400 ;
    END
  END input0[70]
  PIN input0[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 39.6400 75.2400 39.7800 ;
    END
  END input0[69]
  PIN input0[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 34.8300 75.2400 34.9000 ;
    END
  END input0[68]
  PIN input0[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 47.3700 75.2400 47.4400 ;
    END
  END input0[67]
  PIN input0[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT 54.0650 73.9600 54.2050 74.1000 ;
    END
  END input0[66]
  PIN input0[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 52.3850 73.9600 52.5250 74.1000 ;
    END
  END input0[65]
  PIN input0[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 46.4200 74.0300 46.4900 74.1000 ;
    END
  END input0[64]
  PIN input0[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 47.6250 73.9600 47.7650 74.1000 ;
    END
  END input0[63]
  PIN input0[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 42.2400 75.2400 42.3100 ;
    END
  END input0[62]
  PIN input0[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 39.3900 75.2400 39.4600 ;
    END
  END input0[61]
  PIN input0[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 26.2800 74.0300 26.3500 74.1000 ;
    END
  END input0[60]
  PIN input0[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 39.9600 0.0700 40.0300 ;
    END
  END input0[59]
  PIN input0[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 32.2250 73.9600 32.3650 74.1000 ;
    END
  END input0[58]
  PIN input0[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 41.0650 0.1400 41.2050 ;
    END
  END input0[57]
  PIN input0[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 30.0800 75.2400 30.1500 ;
    END
  END input0[56]
  PIN input0[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.5000 0.0000 52.5700 0.0700 ;
    END
  END input0[55]
  PIN input0[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 22.5400 75.2400 22.6800 ;
    END
  END input0[54]
  PIN input0[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 26.2450 75.2400 26.3850 ;
    END
  END input0[53]
  PIN input0[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 33.6550 75.2400 33.7950 ;
    END
  END input0[52]
  PIN input0[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 37.3600 75.2400 37.5000 ;
    END
  END input0[51]
  PIN input0[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 36.9200 74.0300 36.9900 74.1000 ;
    END
  END input0[50]
  PIN input0[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 32.5500 75.2400 32.6200 ;
    END
  END input0[49]
  PIN input0[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 41.1000 75.2400 41.1700 ;
    END
  END input0[48]
  PIN input0[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 49.0800 74.0300 49.1500 74.1000 ;
    END
  END input0[47]
  PIN input0[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 46.9900 74.0300 47.0600 74.1000 ;
    END
  END input0[46]
  PIN input0[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 38.4400 74.0300 38.5100 74.1000 ;
    END
  END input0[45]
  PIN input0[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.3100 74.0300 33.3800 74.1000 ;
    END
  END input0[44]
  PIN input0[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 42.0500 74.0300 42.1200 74.1000 ;
    END
  END input0[43]
  PIN input0[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.2100 74.0300 35.2800 74.1000 ;
    END
  END input0[42]
  PIN input0[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 37.4900 74.0300 37.5600 74.1000 ;
    END
  END input0[41]
  PIN input0[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 38.6300 0.0700 38.7000 ;
    END
  END input0[40]
  PIN input0[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 38.5000 0.1400 38.6400 ;
    END
  END input0[39]
  PIN input0[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.5000 0.0000 33.5700 0.0700 ;
    END
  END input0[38]
  PIN input0[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 36.5400 0.0000 36.6100 0.0700 ;
    END
  END input0[37]
  PIN input0[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 49.8400 0.0000 49.9100 0.0700 ;
    END
  END input0[36]
  PIN input0[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 43.1450 0.0000 43.2850 0.1400 ;
    END
  END input0[35]
  PIN input0[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 45.1050 0.0000 45.2450 0.1400 ;
    END
  END input0[34]
  PIN input0[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 27.4200 75.2400 27.4900 ;
    END
  END input0[33]
  PIN input0[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 29.9500 75.2400 30.0900 ;
    END
  END input0[32]
  PIN input0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 32.5150 75.2400 32.6550 ;
    END
  END input0[31]
  PIN input0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 29.7000 75.2400 29.7700 ;
    END
  END input0[30]
  PIN input0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 36.1600 75.2400 36.2300 ;
    END
  END input0[29]
  PIN input0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 49.4600 74.0300 49.5300 74.1000 ;
    END
  END input0[28]
  PIN input0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 50.9800 75.2400 51.0500 ;
    END
  END input0[27]
  PIN input0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 44.9000 75.2400 44.9700 ;
    END
  END input0[26]
  PIN input0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 46.0400 75.2400 46.1100 ;
    END
  END input0[25]
  PIN input0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 34.2600 74.0300 34.3300 74.1000 ;
    END
  END input0[24]
  PIN input0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 31.4100 74.0300 31.4800 74.1000 ;
    END
  END input0[23]
  PIN input0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 43.1900 74.0300 43.2600 74.1000 ;
    END
  END input0[22]
  PIN input0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 39.9250 0.1400 40.0650 ;
    END
  END input0[21]
  PIN input0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 38.3850 73.9600 38.5250 74.1000 ;
    END
  END input0[20]
  PIN input0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 29.8900 0.0700 29.9600 ;
    END
  END input0[19]
  PIN input0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 29.6650 0.1400 29.8050 ;
    END
  END input0[18]
  PIN input0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 28.7500 0.0700 28.8200 ;
    END
  END input0[17]
  PIN input0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 32.9300 0.0000 33.0000 0.0700 ;
    END
  END input0[16]
  PIN input0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 28.7500 0.0000 28.8200 0.0700 ;
    END
  END input0[15]
  PIN input0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 46.0400 0.0000 46.1100 0.0700 ;
    END
  END input0[14]
  PIN input0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 38.4400 0.0000 38.5100 0.0700 ;
    END
  END input0[13]
  PIN input0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 32.1950 75.2400 32.5950 ;
    END
  END input0[12]
  PIN input0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal9 ;
        RECT 74.4400 32.1850 75.2400 32.9850 ;
    END
  END input0[11]
  PIN input0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 36.2200 75.2400 36.3600 ;
    END
  END input0[10]
  PIN input0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 43.5700 75.2400 43.6400 ;
    END
  END input0[9]
  PIN input0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 42.2050 75.2400 42.3450 ;
    END
  END input0[8]
  PIN input0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 41.0650 75.2400 41.2050 ;
    END
  END input0[7]
  PIN input0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 51.0400 75.2400 51.1800 ;
    END
  END input0[6]
  PIN input0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 45.9100 75.2400 46.0500 ;
    END
  END input0[5]
  PIN input0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.1300 74.0300 48.2000 74.1000 ;
    END
  END input0[4]
  PIN input0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 43.9500 74.0300 44.0200 74.1000 ;
    END
  END input0[3]
  PIN input0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 43.4250 73.9600 43.5650 74.1000 ;
    END
  END input0[2]
  PIN input0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 43.6300 75.2400 43.7700 ;
    END
  END input0[1]
  PIN input0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 38.3850 0.0000 38.5250 0.1400 ;
    END
  END input0[0]
  PIN input1[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 57.8200 0.0700 57.8900 ;
    END
  END input1[79]
  PIN input1[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 62.3800 0.0700 62.4500 ;
    END
  END input1[78]
  PIN input1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 49.6500 0.0700 49.7200 ;
    END
  END input1[77]
  PIN input1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 48.3200 0.0700 48.3900 ;
    END
  END input1[76]
  PIN input1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.0900 0.0000 64.1600 0.0700 ;
    END
  END input1[75]
  PIN input1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 48.5100 0.0000 48.5800 0.0700 ;
    END
  END input1[74]
  PIN input1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 14.1200 75.2400 14.1900 ;
    END
  END input1[73]
  PIN input1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 15.7000 75.2400 15.8400 ;
    END
  END input1[72]
  PIN input1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 29.3450 75.2400 29.7450 ;
    END
  END input1[71]
  PIN input1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 42.6450 75.2400 43.0450 ;
    END
  END input1[70]
  PIN input1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal9 ;
        RECT 74.4400 45.8650 75.2400 46.6650 ;
    END
  END input1[69]
  PIN input1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 38.7850 75.2400 38.9250 ;
    END
  END input1[68]
  PIN input1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 65.6100 74.0300 65.6800 74.1000 ;
    END
  END input1[67]
  PIN input1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 63.9000 75.2400 63.9700 ;
    END
  END input1[66]
  PIN input1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 67.5100 74.0300 67.5800 74.1000 ;
    END
  END input1[65]
  PIN input1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 37.2650 73.9600 37.4050 74.1000 ;
    END
  END input1[64]
  PIN input1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal8 ;
        RECT 47.7750 73.7000 48.1750 74.1000 ;
    END
  END input1[63]
  PIN input1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal9 ;
        RECT 74.4400 42.4450 75.2400 43.2450 ;
    END
  END input1[62]
  PIN input1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 36.3500 0.0700 36.4200 ;
    END
  END input1[61]
  PIN input1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 59.0200 0.1400 59.1600 ;
    END
  END input1[60]
  PIN input1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 47.6200 0.1400 47.7600 ;
    END
  END input1[59]
  PIN input1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 17.3850 73.9600 17.5250 74.1000 ;
    END
  END input1[58]
  PIN input1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 0.0000 57.8450 0.4000 58.2450 ;
    END
  END input1[57]
  PIN input1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 24.2500 75.2400 24.3900 ;
    END
  END input1[56]
  PIN input1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT 60.7850 0.0000 60.9250 0.1400 ;
    END
  END input1[55]
  PIN input1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 11.9950 75.2400 12.1350 ;
    END
  END input1[54]
  PIN input1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 9.4300 75.2400 9.5700 ;
    END
  END input1[53]
  PIN input1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 38.0600 75.2400 38.1300 ;
    END
  END input1[52]
  PIN input1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal9 ;
        RECT 74.4400 37.3150 75.2400 38.1150 ;
    END
  END input1[51]
  PIN input1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 34.2250 0.1400 34.3650 ;
    END
  END input1[50]
  PIN input1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 29.3800 75.2400 29.5200 ;
    END
  END input1[49]
  PIN input1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 45.3400 75.2400 45.4800 ;
    END
  END input1[48]
  PIN input1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 57.9850 73.9600 58.1250 74.1000 ;
    END
  END input1[47]
  PIN input1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal10 ;
        RECT 53.4550 73.3000 54.2550 74.1000 ;
    END
  END input1[46]
  PIN input1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 37.8250 73.9600 37.9650 74.1000 ;
    END
  END input1[45]
  PIN input1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 26.3450 73.9600 26.4850 74.1000 ;
    END
  END input1[44]
  PIN input1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT 47.9050 73.9600 48.0450 74.1000 ;
    END
  END input1[43]
  PIN input1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 29.7050 73.9600 29.8450 74.1000 ;
    END
  END input1[42]
  PIN input1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 29.5100 74.0300 29.5800 74.1000 ;
    END
  END input1[41]
  PIN input1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 0.0000 39.7950 0.4000 40.1950 ;
    END
  END input1[40]
  PIN input1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 35.3650 0.1400 35.5050 ;
    END
  END input1[39]
  PIN input1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 27.1850 0.0000 27.3250 0.1400 ;
    END
  END input1[38]
  PIN input1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 33.3450 0.0000 33.4850 0.1400 ;
    END
  END input1[37]
  PIN input1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 64.4250 0.0000 64.5650 0.1400 ;
    END
  END input1[36]
  PIN input1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 55.7450 0.0000 55.8850 0.1400 ;
    END
  END input1[35]
  PIN input1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 51.8250 0.0000 51.9650 0.1400 ;
    END
  END input1[34]
  PIN input1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 14.5600 75.2400 14.7000 ;
    END
  END input1[33]
  PIN input1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 48.1850 0.0000 48.3250 0.1400 ;
    END
  END input1[32]
  PIN input1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 26.8150 75.2400 26.9550 ;
    END
  END input1[31]
  PIN input1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 27.3850 75.2400 27.5250 ;
    END
  END input1[30]
  PIN input1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal8 ;
        RECT 38.5350 0.0000 38.9350 0.4000 ;
    END
  END input1[29]
  PIN input1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT 58.2650 73.9600 58.4050 74.1000 ;
    END
  END input1[28]
  PIN input1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 66.6650 73.9600 66.8050 74.1000 ;
    END
  END input1[27]
  PIN input1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 53.8900 75.2400 54.0300 ;
    END
  END input1[26]
  PIN input1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 56.4550 75.2400 56.5950 ;
    END
  END input1[25]
  PIN input1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 45.4700 0.0700 45.5400 ;
    END
  END input1[24]
  PIN input1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 26.9050 73.9600 27.0450 74.1000 ;
    END
  END input1[23]
  PIN input1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 42.3050 73.9600 42.4450 74.1000 ;
    END
  END input1[22]
  PIN input1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 28.0250 73.9600 28.1650 74.1000 ;
    END
  END input1[21]
  PIN input1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 36.9850 0.0000 37.1250 0.1400 ;
    END
  END input1[20]
  PIN input1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 23.6200 0.0700 23.6900 ;
    END
  END input1[19]
  PIN input1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 16.2100 0.0700 16.2800 ;
    END
  END input1[18]
  PIN input1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 18.6800 0.0700 18.7500 ;
    END
  END input1[17]
  PIN input1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 23.2400 0.0000 23.3100 0.0700 ;
    END
  END input1[16]
  PIN input1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 16.0200 0.0000 16.0900 0.0700 ;
    END
  END input1[15]
  PIN input1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 51.2650 0.0000 51.4050 0.1400 ;
    END
  END input1[14]
  PIN input1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 37.4900 0.0000 37.5600 0.0700 ;
    END
  END input1[13]
  PIN input1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 29.1300 75.2400 29.2000 ;
    END
  END input1[12]
  PIN input1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 24.8200 75.2400 24.9600 ;
    END
  END input1[11]
  PIN input1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 36.7900 75.2400 36.9300 ;
    END
  END input1[10]
  PIN input1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 41.6350 75.2400 41.7750 ;
    END
  END input1[9]
  PIN input1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 50.1850 75.2400 50.3250 ;
    END
  END input1[8]
  PIN input1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 44.2000 75.2400 44.3400 ;
    END
  END input1[7]
  PIN input1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 57.8450 75.2400 58.2450 ;
    END
  END input1[6]
  PIN input1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal9 ;
        RECT 74.4400 54.4150 75.2400 55.2150 ;
    END
  END input1[5]
  PIN input1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 57.4250 73.9600 57.5650 74.1000 ;
    END
  END input1[4]
  PIN input1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 41.1850 73.9600 41.3250 74.1000 ;
    END
  END input1[3]
  PIN input1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 44.5450 73.9600 44.6850 74.1000 ;
    END
  END input1[2]
  PIN input1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 46.4800 75.2400 46.6200 ;
    END
  END input1[1]
  PIN input1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal6 ;
        RECT 34.1850 0.0000 34.3250 0.1400 ;
    END
  END input1[0]
  PIN ctrl
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 17.4100 0.1400 17.5500 ;
    END
  END ctrl
  PIN output[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 57.4400 0.0700 57.5100 ;
    END
  END output[79]
  PIN output[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 45.0900 0.0700 45.1600 ;
    END
  END output[78]
  PIN output[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 23.4300 74.0300 23.5000 74.1000 ;
    END
  END output[77]
  PIN output[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 50.0300 0.0700 50.1000 ;
    END
  END output[76]
  PIN output[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 18.1100 75.2400 18.1800 ;
    END
  END output[75]
  PIN output[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 70.5500 0.0000 70.6200 0.0700 ;
    END
  END output[74]
  PIN output[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 8.0400 75.2400 8.1100 ;
    END
  END output[73]
  PIN output[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 10.7000 75.2400 10.7700 ;
    END
  END output[72]
  PIN output[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 27.8000 75.2400 27.8700 ;
    END
  END output[71]
  PIN output[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 40.1500 75.2400 40.2200 ;
    END
  END output[70]
  PIN output[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 42.6200 75.2400 42.6900 ;
    END
  END output[69]
  PIN output[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 25.5200 75.2400 25.5900 ;
    END
  END output[68]
  PIN output[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 47.7500 75.2400 47.8200 ;
    END
  END output[67]
  PIN output[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 70.5500 74.0300 70.6200 74.1000 ;
    END
  END output[66]
  PIN output[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 63.3300 74.0300 63.4000 74.1000 ;
    END
  END output[65]
  PIN output[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 51.1700 74.0300 51.2400 74.1000 ;
    END
  END output[64]
  PIN output[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 47.7500 74.0300 47.8200 74.1000 ;
    END
  END output[63]
  PIN output[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.3100 74.0300 52.3800 74.1000 ;
    END
  END output[62]
  PIN output[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 33.6900 74.0300 33.7600 74.1000 ;
    END
  END output[61]
  PIN output[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 25.3300 74.0300 25.4000 74.1000 ;
    END
  END output[60]
  PIN output[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 40.3400 0.0700 40.4100 ;
    END
  END output[59]
  PIN output[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 37.6800 0.0700 37.7500 ;
    END
  END output[58]
  PIN output[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 30.2700 0.0700 30.3400 ;
    END
  END output[57]
  PIN output[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 53.8300 0.0000 53.9000 0.0700 ;
    END
  END output[56]
  PIN output[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 61.0500 0.0000 61.1200 0.0700 ;
    END
  END output[55]
  PIN output[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 70.5850 0.0000 70.7250 0.1400 ;
    END
  END output[54]
  PIN output[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.4100 0.0000 50.4800 0.0700 ;
    END
  END output[53]
  PIN output[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 12.9800 75.2400 13.0500 ;
    END
  END output[52]
  PIN output[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 37.8700 0.0000 37.9400 0.0700 ;
    END
  END output[51]
  PIN output[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 50.7900 0.0000 50.8600 0.0700 ;
    END
  END output[50]
  PIN output[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 43.1900 0.0000 43.2600 0.0700 ;
    END
  END output[49]
  PIN output[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 37.6800 75.2400 37.7500 ;
    END
  END output[48]
  PIN output[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 45.4700 74.0300 45.5400 74.1000 ;
    END
  END output[47]
  PIN output[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 62.5700 74.0300 62.6400 74.1000 ;
    END
  END output[46]
  PIN output[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 54.2100 74.0300 54.2800 74.1000 ;
    END
  END output[45]
  PIN output[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 56.8700 74.0300 56.9400 74.1000 ;
    END
  END output[44]
  PIN output[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 43.5700 74.0300 43.6400 74.1000 ;
    END
  END output[43]
  PIN output[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 28.7500 74.0300 28.8200 74.1000 ;
    END
  END output[42]
  PIN output[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 32.1700 74.0300 32.2400 74.1000 ;
    END
  END output[41]
  PIN output[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 42.6200 0.0700 42.6900 ;
    END
  END output[40]
  PIN output[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 34.0700 0.0000 34.1400 0.0700 ;
    END
  END output[39]
  PIN output[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 30.2700 0.0000 30.3400 0.0700 ;
    END
  END output[38]
  PIN output[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 27.9900 0.0000 28.0600 0.0700 ;
    END
  END output[37]
  PIN output[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 42.4300 0.0000 42.5000 0.0700 ;
    END
  END output[36]
  PIN output[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 45.0900 0.0000 45.1600 0.0700 ;
    END
  END output[35]
  PIN output[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 58.7700 0.0000 58.8400 0.0700 ;
    END
  END output[34]
  PIN output[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 53.4500 0.0000 53.5200 0.0700 ;
    END
  END output[33]
  PIN output[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 41.6700 0.0000 41.7400 0.0700 ;
    END
  END output[32]
  PIN output[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 32.9300 75.2400 33.0000 ;
    END
  END output[31]
  PIN output[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 22.8600 75.2400 22.9300 ;
    END
  END output[30]
  PIN output[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 35.2100 75.2400 35.2800 ;
    END
  END output[29]
  PIN output[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 59.9100 75.2400 59.9800 ;
    END
  END output[28]
  PIN output[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 59.8750 75.2400 60.0150 ;
    END
  END output[27]
  PIN output[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 47.6200 75.2400 47.7600 ;
    END
  END output[26]
  PIN output[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 57.4400 75.2400 57.5100 ;
    END
  END output[25]
  PIN output[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 54.0650 73.9600 54.2050 74.1000 ;
    END
  END output[24]
  PIN output[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 52.6900 74.0300 52.7600 74.1000 ;
    END
  END output[23]
  PIN output[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 45.3850 73.9600 45.5250 74.1000 ;
    END
  END output[22]
  PIN output[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 42.7750 0.1400 42.9150 ;
    END
  END output[21]
  PIN output[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.9700 74.0300 36.0400 74.1000 ;
    END
  END output[20]
  PIN output[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 32.1700 0.0000 32.2400 0.0700 ;
    END
  END output[19]
  PIN output[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 0.0000 30.2350 0.1400 30.3750 ;
    END
  END output[18]
  PIN output[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 22.8600 0.0700 22.9300 ;
    END
  END output[17]
  PIN output[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal4 ;
        RECT 28.0250 0.0000 28.1650 0.1400 ;
    END
  END output[16]
  PIN output[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 0.0000 18.1100 0.0700 18.1800 ;
    END
  END output[15]
  PIN output[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 63.7100 0.0000 63.7800 0.0700 ;
    END
  END output[14]
  PIN output[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 49.2700 0.0000 49.3400 0.0700 ;
    END
  END output[13]
  PIN output[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 17.9800 75.2400 18.1200 ;
    END
  END output[12]
  PIN output[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 15.4500 75.2400 15.5200 ;
    END
  END output[11]
  PIN output[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 27.9550 75.2400 28.0950 ;
    END
  END output[10]
  PIN output[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 42.7750 75.2400 42.9150 ;
    END
  END output[9]
  PIN output[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 47.3950 75.2400 47.7950 ;
    END
  END output[8]
  PIN output[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal5 ;
        RECT 75.1000 40.2100 75.2400 40.3500 ;
    END
  END output[7]
  PIN output[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 59.1500 74.0300 59.2200 74.1000 ;
    END
  END output[6]
  PIN output[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal3 ;
        RECT 75.1700 62.3800 75.2400 62.4500 ;
    END
  END output[5]
  PIN output[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 64.8500 74.0300 64.9200 74.1000 ;
    END
  END output[4]
  PIN output[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 40.1500 74.0300 40.2200 74.1000 ;
    END
  END output[3]
  PIN output[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 45.8500 74.0300 45.9200 74.1000 ;
    END
  END output[2]
  PIN output[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal7 ;
        RECT 74.8400 39.7950 75.2400 40.1950 ;
    END
  END output[1]
  PIN output[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal2 ;
        RECT 35.9700 0.0000 36.0400 0.0700 ;
    END
  END output[0]
  OBS
    LAYER metal10 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal9 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal8 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal7 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal6 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal5 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal4 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal3 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal2 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
    LAYER metal1 ;
      RECT 0.0000 0.0000 75.2400 74.1000 ;
  END
END AsyncMux_width80

END LIBRARY
